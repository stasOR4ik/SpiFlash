`ifndef SPI_FLASH_MEMORY_PKG
`define SPI_FLASH_MEMORY_PKG

package spi_flash_memory_pkg;
	import uvm_pkg::*;

	`include "uvm_macros.svh"

	`include "spi_flash_component.sv"
endpackage

`endif