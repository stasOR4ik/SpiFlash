`ifndef SPI_TRANSACTION
`define SPI_TRANSACTION

class sequence_item;
  byte data;
  time tr_beginning;
endclass;

`endif
